------------------------------------------------------------------------------
--Company:      Loyola Marymount University
--Engineer:     Joseph Gorman

--Create Date:  03/24/2019
--Design Name:
--Module Name:
--Project Name: PCM Communication System
--Tool Versions:
--Description:

--Dependencies:

--Revisions:
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
--use std.textio.all;
--use ieee.std_logic_textio.all;

--entity

--architecture


--open and close file
--architecture test of my_testbench
--  filetest_data_file: text;
--begin
--  file_open(test_data_file, “C:\test.txt”, read_mode);


--assertions will be made to verify transmitted & received data
--assert(transmitted_data) report "It's correct!"
