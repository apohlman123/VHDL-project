------------------------------------------------------------------------------
--Company:      Loyola Marymount University
--Engineer:     Joseph Gorman

--Create Date:  03/24/2019
--Design Name:
--Module Name:
--Project Name: PCM Encoding/Decoding
--Tool Versions:
--Description:

--Dependencies:

--Revisions:
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

--entity

--architecture
